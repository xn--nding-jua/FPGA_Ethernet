-- megafunction wizard: %Triple-Speed Ethernet v13.1%
-- GENERATION: XML
-- PHY_AES50B.vhd

-- Generated using ACDS version 13.1 182 at 2024.12.29.22:38:29

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PHY_AES50B is
	port (
		clk               : in  std_logic                     := '0';             --        control_port_clock_connection.clk
		reset             : in  std_logic                     := '0';             --                     reset_connection.reset
		readdata          : out std_logic_vector(31 downto 0);                    --                         control_port.readdata
		read              : in  std_logic                     := '0';             --                                     .read
		writedata         : in  std_logic_vector(31 downto 0) := (others => '0'); --                                     .writedata
		write             : in  std_logic                     := '0';             --                                     .write
		waitrequest       : out std_logic;                                        --                                     .waitrequest
		address           : in  std_logic_vector(7 downto 0)  := (others => '0'); --                                     .address
		rx_afull_clk      : in  std_logic                     := '0';             -- receive_fifo_status_clock_connection.clk
		rx_afull_data     : in  std_logic_vector(1 downto 0)  := (others => '0'); --                  receive_fifo_status.data
		rx_afull_valid    : in  std_logic                     := '0';             --                                     .valid
		rx_afull_channel  : in  std_logic_vector(0 downto 0)  := (others => '0'); --                                     .channel
		mac_rx_clk_0      : out std_logic;                                        --            mac_rx_clock_connection_0.clk
		mac_tx_clk_0      : out std_logic;                                        --            mac_tx_clock_connection_0.clk
		data_rx_data_0    : out std_logic_vector(7 downto 0);                     --                            receive_0.data
		data_rx_eop_0     : out std_logic;                                        --                                     .endofpacket
		data_rx_error_0   : out std_logic_vector(4 downto 0);                     --                                     .error
		data_rx_ready_0   : in  std_logic                     := '0';             --                                     .ready
		data_rx_sop_0     : out std_logic;                                        --                                     .startofpacket
		data_rx_valid_0   : out std_logic;                                        --                                     .valid
		data_tx_data_0    : in  std_logic_vector(7 downto 0)  := (others => '0'); --                           transmit_0.data
		data_tx_eop_0     : in  std_logic                     := '0';             --                                     .endofpacket
		data_tx_error_0   : in  std_logic                     := '0';             --                                     .error
		data_tx_ready_0   : out std_logic;                                        --                                     .ready
		data_tx_sop_0     : in  std_logic                     := '0';             --                                     .startofpacket
		data_tx_valid_0   : in  std_logic                     := '0';             --                                     .valid
		pkt_class_data_0  : out std_logic_vector(4 downto 0);                     --                receive_packet_type_0.data
		pkt_class_valid_0 : out std_logic;                                        --                                     .valid
		tx_crc_fwd_0      : in  std_logic                     := '0';             --                mac_misc_connection_0.export
		tx_clk_0          : in  std_logic                     := '0';             --        pcs_mac_tx_clock_connection_0.clk
		rx_clk_0          : in  std_logic                     := '0';             --        pcs_mac_rx_clock_connection_0.clk
		set_10_0          : in  std_logic                     := '0';             --              mac_status_connection_0.set_10
		set_1000_0        : in  std_logic                     := '0';             --                                     .set_1000
		eth_mode_0        : out std_logic;                                        --                                     .eth_mode
		ena_10_0          : out std_logic;                                        --                                     .ena_10
		gm_rx_d_0         : in  std_logic_vector(7 downto 0)  := (others => '0'); --                mac_gmii_connection_0.gmii_rx_d
		gm_rx_dv_0        : in  std_logic                     := '0';             --                                     .gmii_rx_dv
		gm_rx_err_0       : in  std_logic                     := '0';             --                                     .gmii_rx_err
		gm_tx_d_0         : out std_logic_vector(7 downto 0);                     --                                     .gmii_tx_d
		gm_tx_en_0        : out std_logic;                                        --                                     .gmii_tx_en
		gm_tx_err_0       : out std_logic;                                        --                                     .gmii_tx_err
		m_rx_d_0          : in  std_logic_vector(3 downto 0)  := (others => '0'); --                 mac_mii_connection_0.mii_rx_d
		m_rx_en_0         : in  std_logic                     := '0';             --                                     .mii_rx_dv
		m_rx_err_0        : in  std_logic                     := '0';             --                                     .mii_rx_err
		m_tx_d_0          : out std_logic_vector(3 downto 0);                     --                                     .mii_tx_d
		m_tx_en_0         : out std_logic;                                        --                                     .mii_tx_en
		m_tx_err_0        : out std_logic;                                        --                                     .mii_tx_err
		mdc               : out std_logic;                                        --                  mac_mdio_connection.mdc
		mdio_in           : in  std_logic                     := '0';             --                                     .mdio_in
		mdio_out          : out std_logic;                                        --                                     .mdio_out
		mdio_oen          : out std_logic                                         --                                     .mdio_oen
	);
end entity PHY_AES50B;

architecture rtl of PHY_AES50B is
	component PHY_AES50B_0002 is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			read              : in  std_logic                     := 'X';             -- read
			writedata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write             : in  std_logic                     := 'X';             -- write
			waitrequest       : out std_logic;                                        -- waitrequest
			address           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			rx_afull_clk      : in  std_logic                     := 'X';             -- clk
			rx_afull_data     : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- data
			rx_afull_valid    : in  std_logic                     := 'X';             -- valid
			rx_afull_channel  : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- channel
			mac_rx_clk_0      : out std_logic;                                        -- clk
			mac_tx_clk_0      : out std_logic;                                        -- clk
			data_rx_data_0    : out std_logic_vector(7 downto 0);                     -- data
			data_rx_eop_0     : out std_logic;                                        -- endofpacket
			data_rx_error_0   : out std_logic_vector(4 downto 0);                     -- error
			data_rx_ready_0   : in  std_logic                     := 'X';             -- ready
			data_rx_sop_0     : out std_logic;                                        -- startofpacket
			data_rx_valid_0   : out std_logic;                                        -- valid
			data_tx_data_0    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			data_tx_eop_0     : in  std_logic                     := 'X';             -- endofpacket
			data_tx_error_0   : in  std_logic                     := 'X';             -- error
			data_tx_ready_0   : out std_logic;                                        -- ready
			data_tx_sop_0     : in  std_logic                     := 'X';             -- startofpacket
			data_tx_valid_0   : in  std_logic                     := 'X';             -- valid
			pkt_class_data_0  : out std_logic_vector(4 downto 0);                     -- data
			pkt_class_valid_0 : out std_logic;                                        -- valid
			tx_crc_fwd_0      : in  std_logic                     := 'X';             -- export
			tx_clk_0          : in  std_logic                     := 'X';             -- clk
			rx_clk_0          : in  std_logic                     := 'X';             -- clk
			set_10_0          : in  std_logic                     := 'X';             -- set_10
			set_1000_0        : in  std_logic                     := 'X';             -- set_1000
			eth_mode_0        : out std_logic;                                        -- eth_mode
			ena_10_0          : out std_logic;                                        -- ena_10
			gm_rx_d_0         : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- gmii_rx_d
			gm_rx_dv_0        : in  std_logic                     := 'X';             -- gmii_rx_dv
			gm_rx_err_0       : in  std_logic                     := 'X';             -- gmii_rx_err
			gm_tx_d_0         : out std_logic_vector(7 downto 0);                     -- gmii_tx_d
			gm_tx_en_0        : out std_logic;                                        -- gmii_tx_en
			gm_tx_err_0       : out std_logic;                                        -- gmii_tx_err
			m_rx_d_0          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_rx_d
			m_rx_en_0         : in  std_logic                     := 'X';             -- mii_rx_dv
			m_rx_err_0        : in  std_logic                     := 'X';             -- mii_rx_err
			m_tx_d_0          : out std_logic_vector(3 downto 0);                     -- mii_tx_d
			m_tx_en_0         : out std_logic;                                        -- mii_tx_en
			m_tx_err_0        : out std_logic;                                        -- mii_tx_err
			mdc               : out std_logic;                                        -- mdc
			mdio_in           : in  std_logic                     := 'X';             -- mdio_in
			mdio_out          : out std_logic;                                        -- mdio_out
			mdio_oen          : out std_logic                                         -- mdio_oen
		);
	end component PHY_AES50B_0002;

begin

	phy_aes50b_inst : component PHY_AES50B_0002
		port map (
			clk               => clk,               --        control_port_clock_connection.clk
			reset             => reset,             --                     reset_connection.reset
			readdata          => readdata,          --                         control_port.readdata
			read              => read,              --                                     .read
			writedata         => writedata,         --                                     .writedata
			write             => write,             --                                     .write
			waitrequest       => waitrequest,       --                                     .waitrequest
			address           => address,           --                                     .address
			rx_afull_clk      => rx_afull_clk,      -- receive_fifo_status_clock_connection.clk
			rx_afull_data     => rx_afull_data,     --                  receive_fifo_status.data
			rx_afull_valid    => rx_afull_valid,    --                                     .valid
			rx_afull_channel  => rx_afull_channel,  --                                     .channel
			mac_rx_clk_0      => mac_rx_clk_0,      --            mac_rx_clock_connection_0.clk
			mac_tx_clk_0      => mac_tx_clk_0,      --            mac_tx_clock_connection_0.clk
			data_rx_data_0    => data_rx_data_0,    --                            receive_0.data
			data_rx_eop_0     => data_rx_eop_0,     --                                     .endofpacket
			data_rx_error_0   => data_rx_error_0,   --                                     .error
			data_rx_ready_0   => data_rx_ready_0,   --                                     .ready
			data_rx_sop_0     => data_rx_sop_0,     --                                     .startofpacket
			data_rx_valid_0   => data_rx_valid_0,   --                                     .valid
			data_tx_data_0    => data_tx_data_0,    --                           transmit_0.data
			data_tx_eop_0     => data_tx_eop_0,     --                                     .endofpacket
			data_tx_error_0   => data_tx_error_0,   --                                     .error
			data_tx_ready_0   => data_tx_ready_0,   --                                     .ready
			data_tx_sop_0     => data_tx_sop_0,     --                                     .startofpacket
			data_tx_valid_0   => data_tx_valid_0,   --                                     .valid
			pkt_class_data_0  => pkt_class_data_0,  --                receive_packet_type_0.data
			pkt_class_valid_0 => pkt_class_valid_0, --                                     .valid
			tx_crc_fwd_0      => tx_crc_fwd_0,      --                mac_misc_connection_0.export
			tx_clk_0          => tx_clk_0,          --        pcs_mac_tx_clock_connection_0.clk
			rx_clk_0          => rx_clk_0,          --        pcs_mac_rx_clock_connection_0.clk
			set_10_0          => set_10_0,          --              mac_status_connection_0.set_10
			set_1000_0        => set_1000_0,        --                                     .set_1000
			eth_mode_0        => eth_mode_0,        --                                     .eth_mode
			ena_10_0          => ena_10_0,          --                                     .ena_10
			gm_rx_d_0         => gm_rx_d_0,         --                mac_gmii_connection_0.gmii_rx_d
			gm_rx_dv_0        => gm_rx_dv_0,        --                                     .gmii_rx_dv
			gm_rx_err_0       => gm_rx_err_0,       --                                     .gmii_rx_err
			gm_tx_d_0         => gm_tx_d_0,         --                                     .gmii_tx_d
			gm_tx_en_0        => gm_tx_en_0,        --                                     .gmii_tx_en
			gm_tx_err_0       => gm_tx_err_0,       --                                     .gmii_tx_err
			m_rx_d_0          => m_rx_d_0,          --                 mac_mii_connection_0.mii_rx_d
			m_rx_en_0         => m_rx_en_0,         --                                     .mii_rx_dv
			m_rx_err_0        => m_rx_err_0,        --                                     .mii_rx_err
			m_tx_d_0          => m_tx_d_0,          --                                     .mii_tx_d
			m_tx_en_0         => m_tx_en_0,         --                                     .mii_tx_en
			m_tx_err_0        => m_tx_err_0,        --                                     .mii_tx_err
			mdc               => mdc,               --                  mac_mdio_connection.mdc
			mdio_in           => mdio_in,           --                                     .mdio_in
			mdio_out          => mdio_out,          --                                     .mdio_out
			mdio_oen          => mdio_oen           --                                     .mdio_oen
		);

end architecture rtl; -- of PHY_AES50B
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2024 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_eth_tse" version="13.1" >
-- Retrieval info: 	<generic name="deviceFamilyName" value="Cyclone III" />
-- Retrieval info: 	<generic name="core_variation" value="MAC_ONLY" />
-- Retrieval info: 	<generic name="ifGMII" value="MII_GMII" />
-- Retrieval info: 	<generic name="enable_use_internal_fifo" value="false" />
-- Retrieval info: 	<generic name="max_channels" value="1" />
-- Retrieval info: 	<generic name="use_misc_ports" value="true" />
-- Retrieval info: 	<generic name="transceiver_type" value="NONE" />
-- Retrieval info: 	<generic name="enable_hd_logic" value="false" />
-- Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
-- Retrieval info: 	<generic name="enable_sup_addr" value="false" />
-- Retrieval info: 	<generic name="stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ext_stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ena_hash" value="false" />
-- Retrieval info: 	<generic name="enable_shift16" value="false" />
-- Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="false" />
-- Retrieval info: 	<generic name="enable_mac_vlan" value="false" />
-- Retrieval info: 	<generic name="enable_magic_detect" value="false" />
-- Retrieval info: 	<generic name="useMDIO" value="true" />
-- Retrieval info: 	<generic name="mdio_clk_div" value="40" />
-- Retrieval info: 	<generic name="enable_ena" value="8" />
-- Retrieval info: 	<generic name="eg_addr" value="11" />
-- Retrieval info: 	<generic name="ing_addr" value="11" />
-- Retrieval info: 	<generic name="phy_identifier" value="0" />
-- Retrieval info: 	<generic name="enable_sgmii" value="false" />
-- Retrieval info: 	<generic name="export_pwrdn" value="false" />
-- Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
-- Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
-- Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
-- Retrieval info: 	<generic name="enable_timestamping" value="false" />
-- Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
-- Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
-- Retrieval info: 	<generic name="AUTO_DEVICE" value="Unknown" />
-- Retrieval info: </instance>
-- IPFS_FILES : PHY_AES50B.vho
-- RELATED_FILES: PHY_AES50B.vhd, PHY_AES50B_0002.v, altera_eth_tse_avalon_arbiter.v, altera_eth_tse_channel_adapter.v, altera_eth_tse_fifoless_mac.v, altera_tse_clk_cntl.v, altera_tse_crc328checker.v, altera_tse_crc328generator.v, altera_tse_crc32ctl8.v, altera_tse_crc32galois8.v, altera_tse_gmii_io.v, altera_tse_lb_read_cntl.v, altera_tse_lb_wrt_cntl.v, altera_tse_hashing.v, altera_tse_host_control.v, altera_tse_host_control_small.v, altera_tse_mac_control.v, altera_tse_register_map.v, altera_tse_register_map_small.v, altera_tse_rx_counter_cntl.v, altera_tse_shared_mac_control.v, altera_tse_shared_register_map.v, altera_tse_tx_counter_cntl.v, altera_tse_lfsr_10.v, altera_tse_loopback_ff.v, altera_tse_altshifttaps.v, altera_tse_fifoless_mac_rx.v, altera_tse_mac_rx.v, altera_tse_fifoless_mac_tx.v, altera_tse_mac_tx.v, altera_tse_magic_detection.v, altera_tse_mdio.v, altera_tse_mdio_clk_gen.v, altera_tse_mdio_cntl.v, altera_tse_top_mdio.v, altera_tse_mii_rx_if.v, altera_tse_mii_tx_if.v, altera_tse_pipeline_base.v, altera_tse_pipeline_stage.sv, altera_tse_dpram_16x32.v, altera_tse_dpram_8x32.v, altera_tse_quad_16x32.v, altera_tse_quad_8x32.v, altera_tse_fifoless_retransmit_cntl.v, altera_tse_retransmit_cntl.v, altera_tse_rgmii_in1.v, altera_tse_rgmii_in4.v, altera_tse_nf_rgmii_module.v, altera_tse_rgmii_module.v, altera_tse_rgmii_out1.v, altera_tse_rgmii_out4.v, altera_tse_rx_ff.v, altera_tse_rx_min_ff.v, altera_tse_rx_ff_cntrl.v, altera_tse_rx_ff_cntrl_32.v, altera_tse_rx_ff_cntrl_32_shift16.v, altera_tse_rx_ff_length.v, altera_tse_rx_stat_extract.v, altera_tse_timing_adapter32.v, altera_tse_timing_adapter8.v, altera_tse_timing_adapter_fifo32.v, altera_tse_timing_adapter_fifo8.v, altera_tse_top_1geth.v, altera_tse_top_fifoless_1geth.v, altera_tse_top_w_fifo.v, altera_tse_top_w_fifo_10_100_1000.v, altera_tse_top_wo_fifo.v, altera_tse_top_wo_fifo_10_100_1000.v, altera_tse_top_gen_host.v, altera_tse_tx_ff.v, altera_tse_tx_min_ff.v, altera_tse_tx_ff_cntrl.v, altera_tse_tx_ff_cntrl_32.v, altera_tse_tx_ff_cntrl_32_shift16.v, altera_tse_tx_ff_length.v, altera_tse_tx_ff_read_cntl.v, altera_tse_tx_stat_extract.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_dc_fifo.v, altera_reset_controller.v, altera_reset_synchronizer.v
